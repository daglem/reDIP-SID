/* verilator lint_off UNUSED */
(* blackbox, keep *)
module SB_WARMBOOT (
	input BOOT,
	input S1,
	input S0
);
endmodule
/* verilator lint_on UNUSED */
